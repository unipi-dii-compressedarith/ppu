module reciprocate_lut #(
        parameter LUT_WIDTH_IN = 8,
        parameter LUT_WIDTH_OUT = 9
    )(
        input [(LUT_WIDTH_IN)-1:0] addr,
        output [(LUT_WIDTH_OUT)-1:0] out   
    );

    reg [(LUT_WIDTH_OUT)-1:0] dout;
    reg [(LUT_WIDTH_OUT)-1:0] mant_recip_rom [(2**LUT_WIDTH_IN - 1):0];

    always @(*) begin 
        case (addr) 
            8'd0 :    dout <= 24'h0;
            8'd1 :    dout <= 24'hff00ff;
            8'd2 :    dout <= 24'hfe03f8;
            8'd3 :    dout <= 24'hfd08e5;
            8'd4 :    dout <= 24'hfc0fc1;
            8'd5 :    dout <= 24'hfb1885;
            8'd6 :    dout <= 24'hfa232d;
            8'd7 :    dout <= 24'hf92fb2;
            8'd8 :    dout <= 24'hf83e10;
            8'd9 :    dout <= 24'hf74e40;
            8'd10 :    dout <= 24'hf6603e;
            8'd11 :    dout <= 24'hf57404;
            8'd12 :    dout <= 24'hf4898d;
            8'd13 :    dout <= 24'hf3a0d5;
            8'd14 :    dout <= 24'hf2b9d6;
            8'd15 :    dout <= 24'hf1d48c;
            8'd16 :    dout <= 24'hf0f0f1;
            8'd17 :    dout <= 24'hf00f01;
            8'd18 :    dout <= 24'hef2eb7;
            8'd19 :    dout <= 24'hee500f;
            8'd20 :    dout <= 24'hed7304;
            8'd21 :    dout <= 24'hec9791;
            8'd22 :    dout <= 24'hebbdb3;
            8'd23 :    dout <= 24'heae564;
            8'd24 :    dout <= 24'hea0ea1;
            8'd25 :    dout <= 24'he93965;
            8'd26 :    dout <= 24'he865ac;
            8'd27 :    dout <= 24'he79373;
            8'd28 :    dout <= 24'he6c2b4;
            8'd29 :    dout <= 24'he5f36d;
            8'd30 :    dout <= 24'he52598;
            8'd31 :    dout <= 24'he45933;
            8'd32 :    dout <= 24'he38e39;
            8'd33 :    dout <= 24'he2c4a7;
            8'd34 :    dout <= 24'he1fc78;
            8'd35 :    dout <= 24'he135aa;
            8'd36 :    dout <= 24'he07038;
            8'd37 :    dout <= 24'hdfac1f;
            8'd38 :    dout <= 24'hdee95c;
            8'd39 :    dout <= 24'hde27eb;
            8'd40 :    dout <= 24'hdd67c9;
            8'd41 :    dout <= 24'hdca8f1;
            8'd42 :    dout <= 24'hdbeb62;
            8'd43 :    dout <= 24'hdb2f17;
            8'd44 :    dout <= 24'hda740e;
            8'd45 :    dout <= 24'hd9ba42;
            8'd46 :    dout <= 24'hd901b2;
            8'd47 :    dout <= 24'hd84a5a;
            8'd48 :    dout <= 24'hd79436;
            8'd49 :    dout <= 24'hd6df44;
            8'd50 :    dout <= 24'hd62b81;
            8'd51 :    dout <= 24'hd578e9;
            8'd52 :    dout <= 24'hd4c77b;
            8'd53 :    dout <= 24'hd41733;
            8'd54 :    dout <= 24'hd3680d;
            8'd55 :    dout <= 24'hd2ba08;
            8'd56 :    dout <= 24'hd20d21;
            8'd57 :    dout <= 24'hd16154;
            8'd58 :    dout <= 24'hd0b6a0;
            8'd59 :    dout <= 24'hd00d01;
            8'd60 :    dout <= 24'hcf6475;
            8'd61 :    dout <= 24'hcebcf9;
            8'd62 :    dout <= 24'hce168a;
            8'd63 :    dout <= 24'hcd7127;
            8'd64 :    dout <= 24'hcccccd;
            8'd65 :    dout <= 24'hcc2978;
            8'd66 :    dout <= 24'hcb8728;
            8'd67 :    dout <= 24'hcae5d8;
            8'd68 :    dout <= 24'hca4588;
            8'd69 :    dout <= 24'hc9a634;
            8'd70 :    dout <= 24'hc907da;
            8'd71 :    dout <= 24'hc86a79;
            8'd72 :    dout <= 24'hc7ce0c;
            8'd73 :    dout <= 24'hc73294;
            8'd74 :    dout <= 24'hc6980c;
            8'd75 :    dout <= 24'hc5fe74;
            8'd76 :    dout <= 24'hc565c8;
            8'd77 :    dout <= 24'hc4ce08;
            8'd78 :    dout <= 24'hc43730;
            8'd79 :    dout <= 24'hc3a13e;
            8'd80 :    dout <= 24'hc30c31;
            8'd81 :    dout <= 24'hc27806;
            8'd82 :    dout <= 24'hc1e4bc;
            8'd83 :    dout <= 24'hc15250;
            8'd84 :    dout <= 24'hc0c0c1;
            8'd85 :    dout <= 24'hc0300c;
            8'd86 :    dout <= 24'hbfa030;
            8'd87 :    dout <= 24'hbf112b;
            8'd88 :    dout <= 24'hbe82fa;
            8'd89 :    dout <= 24'hbdf59d;
            8'd90 :    dout <= 24'hbd6910;
            8'd91 :    dout <= 24'hbcdd53;
            8'd92 :    dout <= 24'hbc5264;
            8'd93 :    dout <= 24'hbbc841;
            8'd94 :    dout <= 24'hbb3ee7;
            8'd95 :    dout <= 24'hbab656;
            8'd96 :    dout <= 24'hba2e8c;
            8'd97 :    dout <= 24'hb9a786;
            8'd98 :    dout <= 24'hb92144;
            8'd99 :    dout <= 24'hb89bc3;
            8'd100 :    dout <= 24'hb81703;
            8'd101 :    dout <= 24'hb79301;
            8'd102 :    dout <= 24'hb70fbb;
            8'd103 :    dout <= 24'hb68d31;
            8'd104 :    dout <= 24'hb60b61;
            8'd105 :    dout <= 24'hb58a48;
            8'd106 :    dout <= 24'hb509e7;
            8'd107 :    dout <= 24'hb48a3a;
            8'd108 :    dout <= 24'hb40b41;
            8'd109 :    dout <= 24'hb38cfa;
            8'd110 :    dout <= 24'hb30f63;
            8'd111 :    dout <= 24'hb2927c;
            8'd112 :    dout <= 24'hb21643;
            8'd113 :    dout <= 24'hb19ab6;
            8'd114 :    dout <= 24'hb11fd4;
            8'd115 :    dout <= 24'hb0a59b;
            8'd116 :    dout <= 24'hb02c0b;
            8'd117 :    dout <= 24'hafb322;
            8'd118 :    dout <= 24'haf3ade;
            8'd119 :    dout <= 24'haec33e;
            8'd120 :    dout <= 24'hae4c41;
            8'd121 :    dout <= 24'hadd5e6;
            8'd122 :    dout <= 24'had602b;
            8'd123 :    dout <= 24'haceb10;
            8'd124 :    dout <= 24'hac7692;
            8'd125 :    dout <= 24'hac02b0;
            8'd126 :    dout <= 24'hab8f6a;
            8'd127 :    dout <= 24'hab1cbe;
            8'd128 :    dout <= 24'haaaaab;
            8'd129 :    dout <= 24'haa392f;
            8'd130 :    dout <= 24'ha9c84a;
            8'd131 :    dout <= 24'ha957fb;
            8'd132 :    dout <= 24'ha8e83f;
            8'd133 :    dout <= 24'ha87917;
            8'd134 :    dout <= 24'ha80a81;
            8'd135 :    dout <= 24'ha79c7b;
            8'd136 :    dout <= 24'ha72f05;
            8'd137 :    dout <= 24'ha6c21e;
            8'd138 :    dout <= 24'ha655c4;
            8'd139 :    dout <= 24'ha5e9f7;
            8'd140 :    dout <= 24'ha57eb5;
            8'd141 :    dout <= 24'ha513fd;
            8'd142 :    dout <= 24'ha4a9cf;
            8'd143 :    dout <= 24'ha44029;
            8'd144 :    dout <= 24'ha3d70a;
            8'd145 :    dout <= 24'ha36e72;
            8'd146 :    dout <= 24'ha3065e;
            8'd147 :    dout <= 24'ha29ecf;
            8'd148 :    dout <= 24'ha237c3;
            8'd149 :    dout <= 24'ha1d13a;
            8'd150 :    dout <= 24'ha16b31;
            8'd151 :    dout <= 24'ha105a9;
            8'd152 :    dout <= 24'ha0a0a1;
            8'd153 :    dout <= 24'ha03c17;
            8'd154 :    dout <= 24'h9fd80a;
            8'd155 :    dout <= 24'h9f747a;
            8'd156 :    dout <= 24'h9f1166;
            8'd157 :    dout <= 24'h9eaecd;
            8'd158 :    dout <= 24'h9e4cad;
            8'd159 :    dout <= 24'h9deb07;
            8'd160 :    dout <= 24'h9d89d9;
            8'd161 :    dout <= 24'h9d2922;
            8'd162 :    dout <= 24'h9cc8e1;
            8'd163 :    dout <= 24'h9c6917;
            8'd164 :    dout <= 24'h9c09c1;
            8'd165 :    dout <= 24'h9baadf;
            8'd166 :    dout <= 24'h9b4c70;
            8'd167 :    dout <= 24'h9aee73;
            8'd168 :    dout <= 24'h9a90e8;
            8'd169 :    dout <= 24'h9a33cd;
            8'd170 :    dout <= 24'h99d723;
            8'd171 :    dout <= 24'h997ae7;
            8'd172 :    dout <= 24'h991f1a;
            8'd173 :    dout <= 24'h98c3bb;
            8'd174 :    dout <= 24'h9868c8;
            8'd175 :    dout <= 24'h980e41;
            8'd176 :    dout <= 24'h97b426;
            8'd177 :    dout <= 24'h975a75;
            8'd178 :    dout <= 24'h97012e;
            8'd179 :    dout <= 24'h96a850;
            8'd180 :    dout <= 24'h964fda;
            8'd181 :    dout <= 24'h95f7cc;
            8'd182 :    dout <= 24'h95a025;
            8'd183 :    dout <= 24'h9548e5;
            8'd184 :    dout <= 24'h94f209;
            8'd185 :    dout <= 24'h949b93;
            8'd186 :    dout <= 24'h944581;
            8'd187 :    dout <= 24'h93efd2;
            8'd188 :    dout <= 24'h939a86;
            8'd189 :    dout <= 24'h93459c;
            8'd190 :    dout <= 24'h92f114;
            8'd191 :    dout <= 24'h929cec;
            8'd192 :    dout <= 24'h924925;
            8'd193 :    dout <= 24'h91f5bd;
            8'd194 :    dout <= 24'h91a2b4;
            8'd195 :    dout <= 24'h915009;
            8'd196 :    dout <= 24'h90fdbc;
            8'd197 :    dout <= 24'h90abcc;
            8'd198 :    dout <= 24'h905a38;
            8'd199 :    dout <= 24'h900901;
            8'd200 :    dout <= 24'h8fb824;
            8'd201 :    dout <= 24'h8f67a2;
            8'd202 :    dout <= 24'h8f177a;
            8'd203 :    dout <= 24'h8ec7ab;
            8'd204 :    dout <= 24'h8e7835;
            8'd205 :    dout <= 24'h8e2918;
            8'd206 :    dout <= 24'h8dda52;
            8'd207 :    dout <= 24'h8d8be3;
            8'd208 :    dout <= 24'h8d3dcb;
            8'd209 :    dout <= 24'h8cf009;
            8'd210 :    dout <= 24'h8ca29c;
            8'd211 :    dout <= 24'h8c5584;
            8'd212 :    dout <= 24'h8c08c1;
            8'd213 :    dout <= 24'h8bbc51;
            8'd214 :    dout <= 24'h8b7034;
            8'd215 :    dout <= 24'h8b246b;
            8'd216 :    dout <= 24'h8ad8f3;
            8'd217 :    dout <= 24'h8a8dcd;
            8'd218 :    dout <= 24'h8a42f8;
            8'd219 :    dout <= 24'h89f874;
            8'd220 :    dout <= 24'h89ae41;
            8'd221 :    dout <= 24'h89645c;
            8'd222 :    dout <= 24'h891ac7;
            8'd223 :    dout <= 24'h88d181;
            8'd224 :    dout <= 24'h888889;
            8'd225 :    dout <= 24'h883fde;
            8'd226 :    dout <= 24'h87f781;
            8'd227 :    dout <= 24'h87af70;
            8'd228 :    dout <= 24'h8767ab;
            8'd229 :    dout <= 24'h872033;
            8'd230 :    dout <= 24'h86d905;
            8'd231 :    dout <= 24'h869223;
            8'd232 :    dout <= 24'h864b8a;
            8'd233 :    dout <= 24'h86053c;
            8'd234 :    dout <= 24'h85bf37;
            8'd235 :    dout <= 24'h85797c;
            8'd236 :    dout <= 24'h853408;
            8'd237 :    dout <= 24'h84eedd;
            8'd238 :    dout <= 24'h84a9fa;
            8'd239 :    dout <= 24'h84655e;
            8'd240 :    dout <= 24'h842108;
            8'd241 :    dout <= 24'h83dcf9;
            8'd242 :    dout <= 24'h839930;
            8'd243 :    dout <= 24'h8355ad;
            8'd244 :    dout <= 24'h83126f;
            8'd245 :    dout <= 24'h82cf75;
            8'd246 :    dout <= 24'h828cc0;
            8'd247 :    dout <= 24'h824a4e;
            8'd248 :    dout <= 24'h820821;
            8'd249 :    dout <= 24'h81c636;
            8'd250 :    dout <= 24'h81848e;
            8'd251 :    dout <= 24'h814328;
            8'd252 :    dout <= 24'h810204;
            8'd253 :    dout <= 24'h80c122;
            8'd254 :    dout <= 24'h808081;
            8'd255 :    dout <= 24'h804020;
            default: 	dout <= 24'h0;
        endcase
    end

    assign out = dout << 1;

endmodule

