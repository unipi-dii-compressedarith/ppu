module fma_posit #(
)(
  input []
);


endmodule: fma_posit
