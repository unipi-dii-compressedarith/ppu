package ppu_pkg;


endpackage