parameter EXP_SIZE_F64 = 11;
parameter MANT_SIZE_F64 = 52;

parameter EXP_SIZE_F32 = 8;
parameter MANT_SIZE_F32 = 23;
