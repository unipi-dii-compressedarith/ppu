/*
Fixed point equivalent values of the rational numbers 
1.466, 1.0012, 2.0 expressed on a range of different bits.

to visualize what i mean try:

>>> import fixed2float as f2f
>>> a = f2f.Fx(3148211028, 1, 32) # e.g.: fp_1_466___N32
>>> print(a, a.eval())


This file exists because SV doesn't support proper conditional compilation.
*/


parameter fp_1_466___N5 = 5'd23;
parameter fp_1_466___N6 = 6'd47;
parameter fp_1_466___N7 = 7'd94;
parameter fp_1_466___N8 = 8'd188;
parameter fp_1_466___N9 = 9'd375;
parameter fp_1_466___N10 = 10'd751;
parameter fp_1_466___N11 = 11'd1501;
parameter fp_1_466___N12 = 12'd3002;
parameter fp_1_466___N13 = 13'd6005;
parameter fp_1_466___N14 = 14'd12009;
parameter fp_1_466___N15 = 15'd24019;
parameter fp_1_466___N16 = 16'd48038;
parameter fp_1_466___N17 = 17'd96076;
parameter fp_1_466___N18 = 18'd192152;
parameter fp_1_466___N19 = 19'd384303;
parameter fp_1_466___N20 = 20'd768606;
parameter fp_1_466___N21 = 21'd1537212;
parameter fp_1_466___N22 = 22'd3074425;
parameter fp_1_466___N23 = 23'd6148850;
parameter fp_1_466___N24 = 24'd12297699;
parameter fp_1_466___N25 = 25'd24595399;
parameter fp_1_466___N26 = 26'd49190797;
parameter fp_1_466___N27 = 27'd98381595;
parameter fp_1_466___N28 = 28'd196763189;
parameter fp_1_466___N29 = 29'd393526378;
parameter fp_1_466___N30 = 30'd787052757;
parameter fp_1_466___N31 = 31'd1574105514;
parameter fp_1_466___N32 = 32'd3148211028;
parameter fp_1_0012___N5 = 9'd256;
parameter fp_1_0012___N6 = 11'd1025;
parameter fp_1_0012___N7 = 13'd4101;
parameter fp_1_0012___N8 = 15'd16404;
parameter fp_1_0012___N9 = 17'd65615;
parameter fp_1_0012___N10 = 19'd262459;
parameter fp_1_0012___N11 = 21'd1049834;
parameter fp_1_0012___N12 = 23'd4199337;
parameter fp_1_0012___N13 = 25'd16797349;
parameter fp_1_0012___N14 = 27'd67189395;
parameter fp_1_0012___N15 = 29'd268757579;
parameter fp_1_0012___N16 = 31'd1075030314;
parameter fp_1_0012___N17 = 33'd4300121257;
parameter fp_1_0012___N18 = 35'd17200485027;
parameter fp_1_0012___N19 = 37'd68801940108;
parameter fp_1_0012___N20 = 39'd275207760432;
parameter fp_1_0012___N21 = 41'd1100831041729;
parameter fp_1_0012___N22 = 43'd4403324166917;
parameter fp_1_0012___N23 = 45'd17613296667669;
parameter fp_1_0012___N24 = 47'd70453186670677;
parameter fp_1_0012___N25 = 49'd281812746682709;
parameter fp_1_0012___N26 = 51'd1127250986730835;
parameter fp_1_0012___N27 = 53'd4509003946923342;
parameter fp_1_0012___N28 = 55'd18036015787693365;
parameter fp_1_0012___N29 = 57'd72144063150773457;
parameter fp_1_0012___N30 = 59'd288576252603093825;
parameter fp_1_0012___N31 = 61'd1154305010412375297;
parameter fp_1_0012___N32 = 63'd4617220041649501185;
parameter fp_2___N5 = 10'd512;
parameter fp_2___N6 = 12'd2048;
parameter fp_2___N7 = 14'd8192;
parameter fp_2___N8 = 16'd32768;
parameter fp_2___N9 = 18'd131072;
parameter fp_2___N10 = 20'd524288;
parameter fp_2___N11 = 22'd2097152;
parameter fp_2___N12 = 24'd8388608;
parameter fp_2___N13 = 26'd33554432;
parameter fp_2___N14 = 28'd134217728;
parameter fp_2___N15 = 30'd536870912;
parameter fp_2___N16 = 32'd2147483648;
parameter fp_2___N17 = 34'd8589934592;
parameter fp_2___N18 = 36'd34359738368;
parameter fp_2___N19 = 38'd137438953472;
parameter fp_2___N20 = 40'd549755813888;
parameter fp_2___N21 = 42'd2199023255552;
parameter fp_2___N22 = 44'd8796093022208;
parameter fp_2___N23 = 46'd35184372088832;
parameter fp_2___N24 = 48'd140737488355328;
parameter fp_2___N25 = 50'd562949953421312;
parameter fp_2___N26 = 52'd2251799813685248;
parameter fp_2___N27 = 54'd9007199254740992;
parameter fp_2___N28 = 56'd36028797018963968;
parameter fp_2___N29 = 58'd144115188075855872;
parameter fp_2___N30 = 60'd576460752303423488;
parameter fp_2___N31 = 62'd2305843009213693952;
parameter fp_2___N32 = 64'd9223372036854775808;
