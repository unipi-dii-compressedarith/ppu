/*

Sat Jan 22 16:55:07 CET 2022

cd waveforms

iverilog -g2012 -DTB_UNSIGNED_RECIPROCAL_APPROX -o unsigned_reciprocal_approx.out \
../src/unsigned_reciprocal_approx.sv \
&& ./unsigned_reciprocal_approx.out

/// WARNING: two numbers are hardcoded and only work in this case with N = 16.

*/



module unsigned_reciprocal_approx #(
        parameter N = 16
    )(
        input [N-1:0] i_data,
        output [N-1:0] o_data
    );

    reg [N-1:0] a, b;
    reg [2*N-1:0] c, d;
    reg [3*N-1:0] e, out;

    assign a = i_data;
    assign b = 16'd48038 - a;
    assign c = $signed(a) * $signed(b);
    assign d = 32'd1075030314 - c;
    assign e = $signed(d) * $signed(b);
    assign out = e << 2;
    
    assign o_data = out[3*N-1: 3*N-1-N];  // (out << 1) >> (2 * N)
endmodule



`ifdef TB_UNSIGNED_RECIPROCAL_APPROX
module tb_unsigned_reciprocal_approx;

    parameter N = 16;

    reg [N-1:0] i_data;
    wire[N-1:0] o_data;


    unsigned_reciprocal_approx unsigned_reciprocal_approx_inst (
        .i_data(i_data),
        .o_data(o_data)
    );


    initial begin
        $dumpfile("tb_unsigned_reciprocal_approx.vcd");
        $dumpvars(0, tb_unsigned_reciprocal_approx);
    end

    // python -c "for i in range(0, 1<<16): print(f\"#10;   i_data = 16'h{hex(i)[2:]};\")" | pbcopy 

    initial begin

  i_data = 16'h0;
#10;   i_data = 16'h1;
#10;   i_data = 16'h4e00;
#10;   i_data = 16'h4e01;
#10;   i_data = 16'h4e02;
#10;   i_data = 16'h4e03;
#10;   i_data = 16'h4e04;
#10;   i_data = 16'h4e05;
#10;   i_data = 16'h4e06;
#10;   i_data = 16'h4e07;
#10;   i_data = 16'h4e08;
#10;   i_data = 16'h4e09;
#10;   i_data = 16'h4e0a;
#10;   i_data = 16'h4e0b;
#10;   i_data = 16'h4e0c;
#10;   i_data = 16'h4e0d;
#10;   i_data = 16'h4e0e;
#10;   i_data = 16'h4e0f;
#10;   i_data = 16'h4e10;
#10;   i_data = 16'h4e11;
#10;   i_data = 16'h4e12;
#10;   i_data = 16'h4e13;
#10;   i_data = 16'h4e14;
#10;   i_data = 16'h4e15;
#10;   i_data = 16'h4e16;
#10;   i_data = 16'h4e17;
#10;   i_data = 16'h4e18;
#10;   i_data = 16'h4e19;
#10;   i_data = 16'h4e1a;
#10;   i_data = 16'h4e1b;
#10;   i_data = 16'h4e1c;
#10;   i_data = 16'h4e1d;
#10;   i_data = 16'h4e1e;
#10;   i_data = 16'h4e1f;
#10;   i_data = 16'h4e20;
#10;   i_data = 16'h4e21;
#10;   i_data = 16'h4e22;
#10;   i_data = 16'h4e23;
#10;   i_data = 16'h4e24;
#10;   i_data = 16'h4e25;
#10;   i_data = 16'h4e26;
#10;   i_data = 16'h4e27;
#10;   i_data = 16'h4e28;
#10;   i_data = 16'h4e29;
#10;   i_data = 16'h4e2a;
#10;   i_data = 16'h4e2b;
#10;   i_data = 16'h4e2c;
#10;   i_data = 16'h4e2d;
#10;   i_data = 16'h4e2e;
#10;   i_data = 16'h4e2f;
#10;   i_data = 16'h4e30;
#10;   i_data = 16'h4e31;
#10;   i_data = 16'h4e32;
#10;   i_data = 16'h4e33;
#10;   i_data = 16'h4e34;
#10;   i_data = 16'h4e35;
#10;   i_data = 16'h4e36;
#10;   i_data = 16'h4e37;
#10;   i_data = 16'h4e38;
#10;   i_data = 16'h4e39;
#10;   i_data = 16'h4e3a;
#10;   i_data = 16'h4e3b;
#10;   i_data = 16'h4e3c;
#10;   i_data = 16'h4e3d;
#10;   i_data = 16'h4e3e;
#10;   i_data = 16'h4e3f;
#10;   i_data = 16'h4e40;
#10;   i_data = 16'h4e41;
#10;   i_data = 16'h4e42;
#10;   i_data = 16'h4e43;
#10;   i_data = 16'h4e44;
#10;   i_data = 16'h4e45;
#10;   i_data = 16'h4e46;
#10;   i_data = 16'h4e47;
#10;   i_data = 16'h4e48;
#10;   i_data = 16'h4e49;
#10;   i_data = 16'h4e4a;
#10;   i_data = 16'h4e4b;
#10;   i_data = 16'h4e4c;
#10;   i_data = 16'h4e4d;
#10;   i_data = 16'h4e4e;
#10;   i_data = 16'h4e4f;
#10;   i_data = 16'h4e50;
#10;   i_data = 16'h4e51;
#10;   i_data = 16'h4e52;
#10;   i_data = 16'h4e53;
#10;   i_data = 16'h4e54;
#10;   i_data = 16'h4e55;
#10;   i_data = 16'h4e56;
#10;   i_data = 16'h4e57;
#10;   i_data = 16'h4e58;
#10;   i_data = 16'h4e59;
#10;   i_data = 16'h4e5a;
#10;   i_data = 16'h4e5b;
#10;   i_data = 16'h4e5c;
#10;   i_data = 16'h4e5d;
#10;   i_data = 16'h4e5e;
#10;   i_data = 16'h4e5f;
#10;   i_data = 16'h4e60;
#10;   i_data = 16'h4e61;
#10;   i_data = 16'h4e62;
#10;   i_data = 16'h4e63;
#10;   i_data = 16'h4e64;
#10;   i_data = 16'h4e65;
#10;   i_data = 16'h4e66;
#10;   i_data = 16'h4e67;
#10;   i_data = 16'h4e68;
#10;   i_data = 16'h4e69;
#10;   i_data = 16'h4e6a;
#10;   i_data = 16'h4e6b;
#10;   i_data = 16'h4e6c;
#10;   i_data = 16'h4e6d;
#10;   i_data = 16'h4e6e;
#10;   i_data = 16'h4e6f;
#10;   i_data = 16'h4e70;
#10;   i_data = 16'h4e71;
#10;   i_data = 16'h4e72;
#10;   i_data = 16'h4e73;
#10;   i_data = 16'h4e74;
#10;   i_data = 16'h4e75;
#10;   i_data = 16'h4e76;
#10;   i_data = 16'h4e77;
#10;   i_data = 16'h4e78;
#10;   i_data = 16'h4e79;
#10;   i_data = 16'h4e7a;
#10;   i_data = 16'h4e7b;
#10;   i_data = 16'h4e7c;
#10;   i_data = 16'h4e7d;
#10;   i_data = 16'h4e7e;
#10;   i_data = 16'h4e7f;
#10;   i_data = 16'h4e80;
#10;   i_data = 16'h4e81;
#10;   i_data = 16'h4e82;
#10;   i_data = 16'h4e83;
#10;   i_data = 16'h4e84;
#10;   i_data = 16'h4e85;
#10;   i_data = 16'h4e86;
#10;   i_data = 16'h4e87;
#10;   i_data = 16'h4e88;
#10;   i_data = 16'h4e89;
#10;   i_data = 16'h4e8a;
#10;   i_data = 16'h4e8b;
#10;   i_data = 16'h4e8c;
#10;   i_data = 16'h4e8d;
#10;   i_data = 16'h4e8e;
#10;   i_data = 16'h4e8f;
#10;   i_data = 16'h4e90;
#10;   i_data = 16'h4e91;
#10;   i_data = 16'h4e92;
#10;   i_data = 16'h4e93;
#10;   i_data = 16'h4e94;
#10;   i_data = 16'h4e95;
#10;   i_data = 16'h4e96;
#10;   i_data = 16'h4e97;
#10;   i_data = 16'h4e98;
#10;   i_data = 16'h4e99;
#10;   i_data = 16'h4e9a;
#10;   i_data = 16'h4e9b;
#10;   i_data = 16'h4e9c;
#10;   i_data = 16'h4e9d;
#10;   i_data = 16'h4e9e;
#10;   i_data = 16'h4e9f;
#10;   i_data = 16'h4ea0;
#10;   i_data = 16'h4ea1;
#10;   i_data = 16'h4ea2;
#10;   i_data = 16'h4ea3;
#10;   i_data = 16'h4ea4;
#10;   i_data = 16'h4ea5;
#10;   i_data = 16'h4ea6;
#10;   i_data = 16'h4ea7;
#10;   i_data = 16'h4ea8;
#10;   i_data = 16'h4ea9;
#10;   i_data = 16'h4eaa;
#10;   i_data = 16'h4eab;
#10;   i_data = 16'h4eac;
#10;   i_data = 16'h4ead;
#10;   i_data = 16'h4eae;
#10;   i_data = 16'h4eaf;
#10;   i_data = 16'h4eb0;
#10;   i_data = 16'h4eb1;
#10;   i_data = 16'h4eb2;
#10;   i_data = 16'h4eb3;
#10;   i_data = 16'h4eb4;
#10;   i_data = 16'h4eb5;
#10;   i_data = 16'h4eb6;
#10;   i_data = 16'h4eb7;
#10;   i_data = 16'h4eb8;
#10;   i_data = 16'h4eb9;
#10;   i_data = 16'h4eba;
#10;   i_data = 16'h4ebb;
#10;   i_data = 16'h4ebc;
#10;   i_data = 16'h4ebd;
#10;   i_data = 16'h4ebe;
#10;   i_data = 16'h4ebf;
#10;   i_data = 16'h4ec0;
#10;   i_data = 16'h4ec1;
#10;   i_data = 16'h4ec2;
#10;   i_data = 16'h4ec3;
#10;   i_data = 16'h4ec4;
#10;   i_data = 16'h4ec5;
#10;   i_data = 16'h4ec6;
#10;   i_data = 16'h4ec7;
#10;   i_data = 16'h4ec8;
#10;   i_data = 16'h4ec9;
#10;   i_data = 16'h4eca;
#10;   i_data = 16'h4ecb;
#10;   i_data = 16'h4ecc;
#10;   i_data = 16'h4ecd;
#10;   i_data = 16'h4ece;
#10;   i_data = 16'h4ecf;
#10;   i_data = 16'h4ed0;
#10;   i_data = 16'h4ed1;
#10;   i_data = 16'h4ed2;
#10;   i_data = 16'h4ed3;
#10;   i_data = 16'h4ed4;
#10;   i_data = 16'h4ed5;
#10;   i_data = 16'h4ed6;
#10;   i_data = 16'h4ed7;
#10;   i_data = 16'h4ed8;
#10;   i_data = 16'h4ed9;
#10;   i_data = 16'h4eda;
#10;   i_data = 16'h4edb;
#10;   i_data = 16'h4edc;
#10;   i_data = 16'h4edd;
#10;   i_data = 16'h4ede;
#10;   i_data = 16'h4edf;
#10;   i_data = 16'h4ee0;
#10;   i_data = 16'h4ee1;
#10;   i_data = 16'h4ee2;
#10;   i_data = 16'h4ee3;
#10;   i_data = 16'h4ee4;
#10;   i_data = 16'h4ee5;
#10;   i_data = 16'h4ee6;
#10;   i_data = 16'h4ee7;
#10;   i_data = 16'h4ee8;
#10;   i_data = 16'h4ee9;
#10;   i_data = 16'h4eea;
#10;   i_data = 16'h4eeb;
#10;   i_data = 16'h4eec;
#10;   i_data = 16'h4eed;
#10;   i_data = 16'h4eee;
#10;   i_data = 16'h4eef;
#10;   i_data = 16'h4ef0;
#10;   i_data = 16'h4ef1;
#10;   i_data = 16'h4ef2;
#10;   i_data = 16'h4ef3;
#10;   i_data = 16'h4ef4;
#10;   i_data = 16'h4ef5;
#10;   i_data = 16'h4ef6;
#10;   i_data = 16'h4ef7;
#10;   i_data = 16'h4ef8;
#10;   i_data = 16'h4ef9;
#10;   i_data = 16'h4efa;
#10;   i_data = 16'h4efb;
#10;   i_data = 16'h4efc;
#10;   i_data = 16'h4efd;
#10;   i_data = 16'h4efe;
#10;   i_data = 16'h4eff;
#10;   i_data = 16'h4f00;
#10;   i_data = 16'h4f01;
#10;   i_data = 16'h4f02;
#10;   i_data = 16'h4f03;
#10;   i_data = 16'h4f04;
#10;   i_data = 16'h4f05;
#10;   i_data = 16'h4f06;
#10;   i_data = 16'h4f07;
#10;   i_data = 16'h4f08;
#10;   i_data = 16'h4f09;
#10;   i_data = 16'h4f0a;
#10;   i_data = 16'h4f0b;
#10;   i_data = 16'h4f0c;
#10;   i_data = 16'h4f0d;
#10;   i_data = 16'h4f0e;
#10;   i_data = 16'h4f0f;
#10;   i_data = 16'h4f10;
#10;   i_data = 16'h4f11;
#10;   i_data = 16'h4f12;
#10;   i_data = 16'h4f13;
#10;   i_data = 16'h4f14;
#10;   i_data = 16'h4f15;
#10;   i_data = 16'h4f16;
#10;   i_data = 16'h4f17;
#10;   i_data = 16'h4f18;
#10;   i_data = 16'h4f19;
#10;   i_data = 16'h4f1a;
#10;   i_data = 16'h4f1b;
#10;   i_data = 16'h4f1c;
#10;   i_data = 16'h4f1d;
#10;   i_data = 16'h4f1e;
#10;   i_data = 16'h4f1f;
#10;   i_data = 16'h4f20;
#10;   i_data = 16'h4f21;
#10;   i_data = 16'h4f22;
#10;   i_data = 16'h4f23;
#10;   i_data = 16'h4f24;
#10;   i_data = 16'h4f25;
#10;   i_data = 16'h4f26;
#10;   i_data = 16'h4f27;
#10;   i_data = 16'h4f28;
#10;   i_data = 16'h4f29;
#10;   i_data = 16'h4f2a;
#10;   i_data = 16'h4f2b;
#10;   i_data = 16'h4f2c;
#10;   i_data = 16'h4f2d;
#10;   i_data = 16'h4f2e;
#10;   i_data = 16'h4f2f;
#10;   i_data = 16'h4f30;
#10;   i_data = 16'h4f31;
#10;   i_data = 16'h4f32;
#10;   i_data = 16'h4f33;
#10;   i_data = 16'h4f34;
#10;   i_data = 16'h4f35;
#10;   i_data = 16'h4f36;
#10;   i_data = 16'h4f37;
#10;   i_data = 16'h4f38;
#10;   i_data = 16'h4f39;
#10;   i_data = 16'h4f3a;
#10;   i_data = 16'h4f3b;
#10;   i_data = 16'h4f3c;
#10;   i_data = 16'h4f3d;
#10;   i_data = 16'h4f3e;
#10;   i_data = 16'h4f3f;
#10;   i_data = 16'h4f40;
#10;   i_data = 16'h4f41;
#10;   i_data = 16'h4f42;
#10;   i_data = 16'h4f43;
#10;   i_data = 16'h4f44;
#10;   i_data = 16'h4f45;
#10;   i_data = 16'h4f46;
#10;   i_data = 16'h4f47;
#10;   i_data = 16'h4f48;
#10;   i_data = 16'h4f49;
#10;   i_data = 16'h4f4a;
#10;   i_data = 16'h4f4b;
#10;   i_data = 16'h4f4c;
#10;   i_data = 16'h4f4d;
#10;   i_data = 16'h4f4e;
#10;   i_data = 16'h4f4f;
#10;   i_data = 16'h4f50;
#10;   i_data = 16'h4f51;
#10;   i_data = 16'h4f52;
#10;   i_data = 16'h4f53;
#10;   i_data = 16'h4f54;
#10;   i_data = 16'h4f55;
#10;   i_data = 16'h4f56;
#10;   i_data = 16'h4f57;
#10;   i_data = 16'h4f58;
#10;   i_data = 16'h4f59;
#10;   i_data = 16'h4f5a;
#10;   i_data = 16'h4f5b;
#10;   i_data = 16'h4f5c;
#10;   i_data = 16'h4f5d;
#10;   i_data = 16'h4f5e;
#10;   i_data = 16'h4f5f;
#10;   i_data = 16'h4f60;
#10;   i_data = 16'h4f61;
#10;   i_data = 16'h4f62;
#10;   i_data = 16'h4f63;
#10;   i_data = 16'h4f64;
#10;   i_data = 16'h4f65;
#10;   i_data = 16'h4f66;
#10;   i_data = 16'h4f67;
#10;   i_data = 16'h4f68;
#10;   i_data = 16'h4f69;
#10;   i_data = 16'h4f6a;
#10;   i_data = 16'h4f6b;
#10;   i_data = 16'h4f6c;
#10;   i_data = 16'h4f6d;
#10;   i_data = 16'h4f6e;
#10;   i_data = 16'h4f6f;
#10;   i_data = 16'h4f70;
#10;   i_data = 16'h4f71;
#10;   i_data = 16'h4f72;
#10;   i_data = 16'h4f73;
#10;   i_data = 16'h4f74;
#10;   i_data = 16'h4f75;
#10;   i_data = 16'h4f76;
#10;   i_data = 16'h4f77;
#10;   i_data = 16'h4f78;
#10;   i_data = 16'h4f79;
#10;   i_data = 16'h4f7a;
#10;   i_data = 16'h4f7b;
#10;   i_data = 16'h4f7c;
#10;   i_data = 16'h4f7d;
#10;   i_data = 16'h4f7e;
#10;   i_data = 16'h4f7f;
#10;   i_data = 16'h4f80;
#10;   i_data = 16'h4f81;
#10;   i_data = 16'h4f82;
#10;   i_data = 16'h4f83;
#10;   i_data = 16'h4f84;
#10;   i_data = 16'h4f85;
#10;   i_data = 16'h4f86;
#10;   i_data = 16'h4f87;
#10;   i_data = 16'h4f88;
#10;   i_data = 16'h4f89;
#10;   i_data = 16'h4f8a;
#10;   i_data = 16'h4f8b;
#10;   i_data = 16'h4f8c;
#10;   i_data = 16'h4f8d;
#10;   i_data = 16'h4f8e;
#10;   i_data = 16'h4f8f;
#10;   i_data = 16'h4f90;
#10;   i_data = 16'h4f91;
#10;   i_data = 16'h4f92;
#10;   i_data = 16'h4f93;
#10;   i_data = 16'h4f94;
#10;   i_data = 16'h4f95;
#10;   i_data = 16'h4f96;
#10;   i_data = 16'h4f97;
#10;   i_data = 16'h4f98;
#10;   i_data = 16'h4f99;
#10;   i_data = 16'h4f9a;
#10;   i_data = 16'h4f9b;
#10;   i_data = 16'h4f9c;
#10;   i_data = 16'h4f9d;
#10;   i_data = 16'h4f9e;
#10;   i_data = 16'h4f9f;
#10;   i_data = 16'h4fa0;
#10;   i_data = 16'h4fa1;
#10;   i_data = 16'h4fa2;
#10;   i_data = 16'h4fa3;
#10;   i_data = 16'h4fa4;
#10;   i_data = 16'h4fa5;
#10;   i_data = 16'h4fa6;
#10;   i_data = 16'h4fa7;
#10;   i_data = 16'h4fa8;
#10;   i_data = 16'h4fa9;
#10;   i_data = 16'h4faa;
#10;   i_data = 16'h4fab;
#10;   i_data = 16'h4fac;
#10;   i_data = 16'h4fad;
#10;   i_data = 16'h4fae;
#10;   i_data = 16'h4faf;
#10;   i_data = 16'h4fb0;
#10;   i_data = 16'h4fb1;
#10;   i_data = 16'h4fb2;
#10;   i_data = 16'h4fb3;
#10;   i_data = 16'h4fb4;
#10;   i_data = 16'h4fb5;
#10;   i_data = 16'h4fb6;
#10;   i_data = 16'h4fb7;
#10;   i_data = 16'h4fb8;
#10;   i_data = 16'h4fb9;
#10;   i_data = 16'h4fba;
#10;   i_data = 16'h4fbb;
#10;   i_data = 16'h4fbc;
#10;   i_data = 16'h4fbd;
#10;   i_data = 16'h4fbe;
#10;   i_data = 16'h4fbf;
#10;   i_data = 16'h4fc0;
#10;   i_data = 16'h4fc1;
#10;   i_data = 16'h4fc2;
#10;   i_data = 16'h4fc3;
#10;   i_data = 16'h4fc4;
#10;   i_data = 16'h4fc5;
#10;   i_data = 16'h4fc6;
#10;   i_data = 16'h4fc7;
#10;   i_data = 16'h4fc8;
#10;   i_data = 16'h4fc9;
#10;   i_data = 16'h4fca;
#10;   i_data = 16'h4fcb;
#10;   i_data = 16'h4fcc;
#10;   i_data = 16'h4fcd;
#10;   i_data = 16'h4fce;
#10;   i_data = 16'h4fcf;
#10;   i_data = 16'h4fd0;
#10;   i_data = 16'h4fd1;
#10;   i_data = 16'h4fd2;
#10;   i_data = 16'h4fd3;
#10;   i_data = 16'h4fd4;
#10;   i_data = 16'h4fd5;
#10;   i_data = 16'h4fd6;
#10;   i_data = 16'h4fd7;
#10;   i_data = 16'h4fd8;
#10;   i_data = 16'h4fd9;
#10;   i_data = 16'h4fda;
#10;   i_data = 16'h4fdb;
#10;   i_data = 16'h4fdc;
#10;   i_data = 16'h4fdd;
#10;   i_data = 16'h4fde;
#10;   i_data = 16'h4fdf;
#10;   i_data = 16'h4fe0;
#10;   i_data = 16'h4fe1;
#10;   i_data = 16'h4fe2;
#10;   i_data = 16'h4fe3;
#10;   i_data = 16'h4fe4;
#10;   i_data = 16'h4fe5;
#10;   i_data = 16'h4fe6;
#10;   i_data = 16'h4fe7;
#10;   i_data = 16'h4fe8;
#10;   i_data = 16'h4fe9;
#10;   i_data = 16'h4fea;
#10;   i_data = 16'h4feb;
#10;   i_data = 16'h4fec;
#10;   i_data = 16'h4fed;
#10;   i_data = 16'h4fee;
#10;   i_data = 16'h4fef;
#10;   i_data = 16'h4ff0;
#10;   i_data = 16'h4ff1;
#10;   i_data = 16'h4ff2;
#10;   i_data = 16'h4ff3;
#10;   i_data = 16'h4ff4;
#10;   i_data = 16'h4ff5;
#10;   i_data = 16'h4ff6;
#10;   i_data = 16'h4ff7;
#10;   i_data = 16'h4ff8;
#10;   i_data = 16'h4ff9;
#10;   i_data = 16'h4ffa;
#10;   i_data = 16'h4ffb;
#10;   i_data = 16'h4ffc;
#10;   i_data = 16'h4ffd;
#10;   i_data = 16'h4ffe;
#10;   i_data = 16'h4fff;
#10;   i_data = 16'h5000;
#10;   i_data = 16'h5001;
#10;   i_data = 16'h5002;
#10;   i_data = 16'h5003;
#10;   i_data = 16'h5004;
#10;   i_data = 16'h5005;
#10;   i_data = 16'h5006;
#10;   i_data = 16'h5007;
#10;   i_data = 16'h5008;
#10;   i_data = 16'h5009;
#10;   i_data = 16'h500a;
#10;   i_data = 16'h500b;
#10;   i_data = 16'h500c;
#10;   i_data = 16'h500d;
#10;   i_data = 16'h500e;
#10;   i_data = 16'h500f;
#10;   i_data = 16'h5010;
#10;   i_data = 16'h5011;
#10;   i_data = 16'h5012;
#10;   i_data = 16'h5013;
#10;   i_data = 16'h5014;
#10;   i_data = 16'h5015;
#10;   i_data = 16'h5016;
#10;   i_data = 16'h5017;
#10;   i_data = 16'h5018;
#10;   i_data = 16'h5019;
#10;   i_data = 16'h501a;
#10;   i_data = 16'h501b;
#10;   i_data = 16'h501c;
#10;   i_data = 16'h501d;
#10;   i_data = 16'h501e;
#10;   i_data = 16'h501f;
#10;   i_data = 16'h5020;
#10;   i_data = 16'h5021;
#10;   i_data = 16'h5022;
#10;   i_data = 16'h5023;
#10;   i_data = 16'h5024;
#10;   i_data = 16'h5025;
#10;   i_data = 16'h5026;
#10;   i_data = 16'h5027;
#10;   i_data = 16'h5028;
#10;   i_data = 16'h5029;
#10;   i_data = 16'h502a;
#10;   i_data = 16'h502b;
#10;   i_data = 16'h502c;
#10;   i_data = 16'h502d;
#10;   i_data = 16'h502e;
#10;   i_data = 16'h502f;
#10;   i_data = 16'h5030;
#10;   i_data = 16'h5031;
#10;   i_data = 16'h5032;
#10;   i_data = 16'h5033;
#10;   i_data = 16'h5034;
#10;   i_data = 16'h5035;
#10;   i_data = 16'h5036;
#10;   i_data = 16'h5037;
#10;   i_data = 16'h5038;
#10;   i_data = 16'h5039;
#10;   i_data = 16'h503a;
#10;   i_data = 16'h503b;
#10;   i_data = 16'h503c;
#10;   i_data = 16'h503d;
#10;   i_data = 16'h503e;
#10;   i_data = 16'h503f;
#10;   i_data = 16'h5040;
#10;   i_data = 16'h5041;
#10;   i_data = 16'h5042;
#10;   i_data = 16'h5043;
#10;   i_data = 16'h5044;
#10;   i_data = 16'h5045;
#10;   i_data = 16'h5046;
#10;   i_data = 16'h5047;
#10;   i_data = 16'h5048;
#10;   i_data = 16'h5049;
#10;   i_data = 16'h504a;
#10;   i_data = 16'h504b;
#10;   i_data = 16'h504c;
#10;   i_data = 16'h504d;
#10;   i_data = 16'h504e;
#10;   i_data = 16'h504f;
#10;   i_data = 16'h5050;
#10;   i_data = 16'h5051;
#10;   i_data = 16'h5052;
#10;   i_data = 16'h5053;
#10;   i_data = 16'h5054;
#10;   i_data = 16'h5055;
#10;   i_data = 16'h5056;
#10;   i_data = 16'h5057;
#10;   i_data = 16'h5058;
#10;   i_data = 16'h5059;
#10;   i_data = 16'h505a;
#10;   i_data = 16'h505b;
#10;   i_data = 16'h505c;
#10;   i_data = 16'h505d;
#10;   i_data = 16'h505e;
#10;   i_data = 16'h505f;
#10;   i_data = 16'h5060;
#10;   i_data = 16'h5061;
#10;   i_data = 16'h5062;
#10;   i_data = 16'h5063;
#10;   i_data = 16'h5064;
#10;   i_data = 16'h5065;
#10;   i_data = 16'h5066;
#10;   i_data = 16'h5067;
#10;   i_data = 16'h5068;
#10;   i_data = 16'h5069;
#10;   i_data = 16'h506a;
#10;   i_data = 16'h506b;
#10;   i_data = 16'h506c;
#10;   i_data = 16'h506d;
#10;   i_data = 16'h506e;
#10;   i_data = 16'h506f;
#10;   i_data = 16'h5070;
#10;   i_data = 16'h5071;
#10;   i_data = 16'h5072;
#10;   i_data = 16'h5073;
#10;   i_data = 16'h5074;
#10;   i_data = 16'h5075;
#10;   i_data = 16'h5076;
#10;   i_data = 16'h5077;
#10;   i_data = 16'h5078;
#10;   i_data = 16'h5079;
#10;   i_data = 16'h507a;
#10;   i_data = 16'h507b;
#10;   i_data = 16'h507c;
#10;   i_data = 16'h507d;
#10;   i_data = 16'h507e;
#10;   i_data = 16'h507f;
#10;   i_data = 16'h5080;
#10;   i_data = 16'h5081;
#10;   i_data = 16'h5082;
#10;   i_data = 16'h5083;
#10;   i_data = 16'h5084;
#10;   i_data = 16'h5085;
#10;   i_data = 16'h5086;
#10;   i_data = 16'h5087;
#10;   i_data = 16'h5088;
#10;   i_data = 16'h5089;
#10;   i_data = 16'h508a;
#10;   i_data = 16'h508b;
#10;   i_data = 16'h508c;
#10;   i_data = 16'h508d;
#10;   i_data = 16'h508e;
#10;   i_data = 16'h508f;
#10;   i_data = 16'h5090;
#10;   i_data = 16'h5091;
#10;   i_data = 16'h5092;
#10;   i_data = 16'h5093;
#10;   i_data = 16'h5094;
#10;   i_data = 16'h5095;
#10;   i_data = 16'h5096;
#10;   i_data = 16'h5097;
#10;   i_data = 16'h5098;
#10;   i_data = 16'h5099;
#10;   i_data = 16'h509a;
#10;   i_data = 16'h509b;
#10;   i_data = 16'h509c;
#10;   i_data = 16'h509d;
#10;   i_data = 16'h509e;
#10;   i_data = 16'h509f;
#10;   i_data = 16'h50a0;
#10;   i_data = 16'h50a1;
#10;   i_data = 16'h50a2;
#10;   i_data = 16'h50a3;
#10;   i_data = 16'h50a4;
#10;   i_data = 16'h50a5;
#10;   i_data = 16'h50a6;
#10;   i_data = 16'h50a7;
#10;   i_data = 16'h50a8;
#10;   i_data = 16'h50a9;
#10;   i_data = 16'h50aa;
#10;   i_data = 16'h50ab;
#10;   i_data = 16'h50ac;
#10;   i_data = 16'h50ad;
#10;   i_data = 16'h50ae;
#10;   i_data = 16'h50af;
#10;   i_data = 16'h50b0;
#10;   i_data = 16'h50b1;
#10;   i_data = 16'h50b2;
#10;   i_data = 16'h50b3;
#10;   i_data = 16'h50b4;
#10;   i_data = 16'h50b5;
#10;   i_data = 16'h50b6;
#10;   i_data = 16'h50b7;
#10;   i_data = 16'h50b8;
#10;   i_data = 16'h50b9;
#10;   i_data = 16'h50ba;
#10;   i_data = 16'h50bb;
#10;   i_data = 16'h50bc;
#10;   i_data = 16'h50bd;
#10;   i_data = 16'h50be;
#10;   i_data = 16'h50bf;
#10;   i_data = 16'h50c0;
#10;   i_data = 16'h50c1;
#10;   i_data = 16'h50c2;
#10;   i_data = 16'h50c3;
#10;   i_data = 16'h50c4;
#10;   i_data = 16'h50c5;
#10;   i_data = 16'h50c6;
#10;   i_data = 16'h50c7;
#10;   i_data = 16'h50c8;
#10;   i_data = 16'h50c9;
#10;   i_data = 16'h50ca;
#10;   i_data = 16'h50cb;
#10;   i_data = 16'h50cc;
#10;   i_data = 16'h50cd;
#10;   i_data = 16'h50ce;
#10;   i_data = 16'h50cf;
#10;   i_data = 16'h50d0;
#10;   i_data = 16'h50d1;
#10;   i_data = 16'h50d2;
#10;   i_data = 16'h50d3;
#10;   i_data = 16'h50d4;
#10;   i_data = 16'h50d5;
#10;   i_data = 16'h50d6;
#10;   i_data = 16'h50d7;
#10;   i_data = 16'h50d8;
#10;   i_data = 16'h50d9;
#10;   i_data = 16'h50da;
#10;   i_data = 16'h50db;
#10;   i_data = 16'h50dc;
#10;   i_data = 16'h50dd;
#10;   i_data = 16'h50de;
#10;   i_data = 16'h50df;
#10;   i_data = 16'h50e0;
#10;   i_data = 16'h50e1;
#10;   i_data = 16'h50e2;
#10;   i_data = 16'h50e3;
#10;   i_data = 16'h50e4;
#10;   i_data = 16'h50e5;
#10;   i_data = 16'h50e6;
#10;   i_data = 16'h50e7;
#10;   i_data = 16'h50e8;
#10;   i_data = 16'h50e9;
#10;   i_data = 16'h50ea;
#10;   i_data = 16'h50eb;
#10;   i_data = 16'h50ec;
#10;   i_data = 16'h50ed;
#10;   i_data = 16'h50ee;
#10;   i_data = 16'h50ef;
#10;   i_data = 16'h50f0;
#10;   i_data = 16'h50f1;
#10;   i_data = 16'h50f2;
#10;   i_data = 16'h50f3;
#10;   i_data = 16'h50f4;
#10;   i_data = 16'h50f5;
#10;   i_data = 16'h50f6;
#10;   i_data = 16'h50f7;
#10;   i_data = 16'h50f8;
#10;   i_data = 16'h50f9;
#10;   i_data = 16'h50fa;
#10;   i_data = 16'h50fb;
#10;   i_data = 16'h50fc;
#10;   i_data = 16'h50fd;
#10;   i_data = 16'h50fe;
#10;   i_data = 16'h50ff;
#10;   i_data = 16'h5100;
#10;   i_data = 16'h5101;
#10;   i_data = 16'h5102;
#10;   i_data = 16'h5103;
#10;   i_data = 16'h5104;
#10;   i_data = 16'h5105;
#10;   i_data = 16'h5106;
#10;   i_data = 16'h5107;
#10;   i_data = 16'h5108;
#10;   i_data = 16'h5109;
#10;   i_data = 16'h510a;
#10;   i_data = 16'h510b;
#10;   i_data = 16'h510c;
#10;   i_data = 16'h510d;
#10;   i_data = 16'h510e;
#10;   i_data = 16'h510f;
#10;   i_data = 16'h5110;
#10;   i_data = 16'h5111;
#10;   i_data = 16'h5112;
#10;   i_data = 16'h5113;
#10;   i_data = 16'h5114;
#10;   i_data = 16'h5115;
#10;   i_data = 16'h5116;
#10;   i_data = 16'h5117;
#10;   i_data = 16'h5118;
#10;   i_data = 16'h5119;
#10;   i_data = 16'h511a;
#10;   i_data = 16'h511b;
#10;   i_data = 16'h511c;
#10;   i_data = 16'h511d;
#10;   i_data = 16'h511e;
#10;   i_data = 16'h511f;
#10;   i_data = 16'h5120;
#10;   i_data = 16'h5121;
#10;   i_data = 16'h5122;
#10;   i_data = 16'h5123;
#10;   i_data = 16'h5124;
#10;   i_data = 16'h5125;
#10;   i_data = 16'h5126;
#10;   i_data = 16'h5127;
#10;   i_data = 16'h5128;
#10;   i_data = 16'h5129;
#10;   i_data = 16'h512a;
#10;   i_data = 16'h512b;
#10;   i_data = 16'h512c;
#10;   i_data = 16'h512d;
#10;   i_data = 16'h512e;
#10;   i_data = 16'h512f;
#10;   i_data = 16'h5130;
#10;   i_data = 16'h5131;
#10;   i_data = 16'h5132;
#10;   i_data = 16'h5133;
#10;   i_data = 16'h5134;
#10;   i_data = 16'h5135;
#10;   i_data = 16'h5136;
#10;   i_data = 16'h5137;
#10;   i_data = 16'h5138;
#10;   i_data = 16'h5139;
#10;   i_data = 16'h513a;
#10;   i_data = 16'h513b;
#10;   i_data = 16'h513c;
#10;
end

endmodule
`endif
