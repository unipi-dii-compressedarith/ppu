/*
Fixed point equivalent values of the rational numbers
1.466, 1.0012, 2.0 expressed on a range of different bits.

to visualize what i mean try:

>>> import fixed2float as f2f
>>> a = f2f.Fx(3148211028, 1, 32) # e.g.: fx_1_466___N32
>>> print(a, a.eval())


This file exists because SV doesn't support proper conditional compilation.
*/






parameter fx_1_466___N5 = 3'd6;
parameter fx_1_466___N6 = 4'd12;
parameter fx_1_466___N7 = 5'd23;
parameter fx_1_466___N8 = 6'd47;
parameter fx_1_466___N9 = 7'd94;
parameter fx_1_466___N10 = 8'd188;
parameter fx_1_466___N11 = 9'd375;
parameter fx_1_466___N12 = 10'd751;
parameter fx_1_466___N13 = 11'd1501;
parameter fx_1_466___N14 = 12'd3002;
parameter fx_1_466___N15 = 13'd6005;
parameter fx_1_466___N16 = 14'd12009;
parameter fx_1_466___N17 = 15'd24019;
parameter fx_1_466___N18 = 16'd48038;
parameter fx_1_466___N19 = 17'd96076;
parameter fx_1_466___N20 = 18'd192152;
parameter fx_1_466___N21 = 19'd384303;
parameter fx_1_466___N22 = 20'd768606;
parameter fx_1_466___N23 = 21'd1537212;
parameter fx_1_466___N24 = 22'd3074425;
parameter fx_1_466___N25 = 23'd6148850;
parameter fx_1_466___N26 = 24'd12297699;
parameter fx_1_466___N27 = 25'd24595399;
parameter fx_1_466___N28 = 26'd49190797;
parameter fx_1_466___N29 = 27'd98381595;
parameter fx_1_466___N30 = 28'd196763189;
parameter fx_1_466___N31 = 29'd393526378;
parameter fx_1_466___N32 = 30'd787052757;

parameter fx_1_0012___N5 = 5'd16;
parameter fx_1_0012___N6 = 7'd64;
parameter fx_1_0012___N7 = 9'd256;
parameter fx_1_0012___N8 = 11'd1025;
parameter fx_1_0012___N9 = 13'd4101;
parameter fx_1_0012___N10 = 15'd16404;
parameter fx_1_0012___N11 = 17'd65615;
parameter fx_1_0012___N12 = 19'd262459;
parameter fx_1_0012___N13 = 21'd1049834;
parameter fx_1_0012___N14 = 23'd4199337;
parameter fx_1_0012___N15 = 25'd16797349;
parameter fx_1_0012___N16 = 27'd67189395;
parameter fx_1_0012___N17 = 29'd268757579;
parameter fx_1_0012___N18 = 31'd1075030314;
parameter fx_1_0012___N19 = 33'd4300121257;
parameter fx_1_0012___N20 = 35'd17200485027;
parameter fx_1_0012___N21 = 37'd68801940108;
parameter fx_1_0012___N22 = 39'd275207760432;
parameter fx_1_0012___N23 = 41'd1100831041729;
parameter fx_1_0012___N24 = 43'd4403324166917;
parameter fx_1_0012___N25 = 45'd17613296667669;
parameter fx_1_0012___N26 = 47'd70453186670677;
parameter fx_1_0012___N27 = 49'd281812746682709;
parameter fx_1_0012___N28 = 51'd1127250986730835;
parameter fx_1_0012___N29 = 53'd4509003946923342;
parameter fx_1_0012___N30 = 55'd18036015787693365;
parameter fx_1_0012___N31 = 57'd72144063150773457;
parameter fx_1_0012___N32 = 59'd288576252603093825;

parameter fx_2___N5 = 6'd32;
parameter fx_2___N6 = 8'd128;
parameter fx_2___N7 = 10'd512;
parameter fx_2___N8 = 12'd2048;
parameter fx_2___N9 = 14'd8192;
parameter fx_2___N10 = 16'd32768;
parameter fx_2___N11 = 18'd131072;
parameter fx_2___N12 = 20'd524288;
parameter fx_2___N13 = 22'd2097152;
parameter fx_2___N14 = 24'd8388608;
parameter fx_2___N15 = 26'd33554432;
parameter fx_2___N16 = 28'd134217728;
parameter fx_2___N17 = 30'd536870912;
parameter fx_2___N18 = 32'd2147483648;
parameter fx_2___N19 = 34'd8589934592;
parameter fx_2___N20 = 36'd34359738368;
parameter fx_2___N21 = 38'd137438953472;
parameter fx_2___N22 = 40'd549755813888;
parameter fx_2___N23 = 42'd2199023255552;
parameter fx_2___N24 = 44'd8796093022208;
parameter fx_2___N25 = 46'd35184372088832;
parameter fx_2___N26 = 48'd140737488355328;
parameter fx_2___N27 = 50'd562949953421312;
parameter fx_2___N28 = 52'd2251799813685248;
parameter fx_2___N29 = 54'd9007199254740992;
parameter fx_2___N30 = 56'd36028797018963968;
parameter fx_2___N31 = 58'd144115188075855872;
parameter fx_2___N32 = 60'd576460752303423488;
