import p8e0_pkg::*;

module p8e0_add(
        input        [7:0]    a,
        input        [7:0]    b,
        output /* wire */     is_zero,
        output    wire        is_nar,
        output logic [7:0]    z
    );






endmodule