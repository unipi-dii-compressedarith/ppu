parameter FLOAT_EXP_SIZE_F64 = 11;
parameter FLOAT_MANT_SIZE_F64 = 52;

parameter FLOAT_EXP_SIZE_F32 = 8;
parameter FLOAT_MANT_SIZE_F32 = 23;

parameter FLOAT_EXP_SIZE_F16 = 5;
parameter FLOAT_MANT_SIZE_F16 = 10;
