module core_sub #(
        parameter N = 4
    )(
        input [(MANT_ADD_RESULT_SIZE-1)-1:0] mant,
        input [TE_SIZE-1:0] te_diff,
        output [(MANT_ADD_RESULT_SIZE)-1:0] new_mant,
        output [TE_SIZE-1:0] new_te_diff
    );

    wire [($clog2(MANT_ADD_RESULT_SIZE-1))-1:0] leading_zeros;

    cls #(
        .NUM_BITS(MANT_ADD_RESULT_SIZE-1)
    ) clz (
        .bits               (mant),
        .val                (1'b0),
        .leading_set        (leading_zeros),
        .index_highest_set  ()
    );

    assign new_te_diff = te_diff - leading_zeros;
    assign new_mant = (mant << leading_zeros); // & ~(1 << (MANT_SUB_RESULT_SIZE-1));

endmodule
